`timescale 1ns / 100ps
`default_nettype none

module fmv_w_s (x, y);
    input wire [31:0] x;
    output [31:0] y;

    wire [31:0] y;

    assign y = x;
endmodule
